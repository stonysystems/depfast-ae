#include<__dep__.h>
#include "eRPC"
class ExampleClientServiceImplWrapper{

    ExampleClientServiceImplWrapper()
    void hello(const std::vector<int32_t>& _req, erpc::ReqHandle *req_handle)    
};